module encoder {
	
};
endmodule